module level_4(
    input [63:0] temp_3, output [63:0] temp_4
);

    parallel_prefix mod96(temp_3[3:2], 2'b00, temp_4[3:2]);
    parallel_prefix mod97(temp_3[3:2], 2'b00, temp_4[3:2]);
    parallel_prefix mod98(temp_3[5:4], 2'b00, temp_4[5:4]);
    parallel_prefix mod99(temp_3[7:6], 2'b00, temp_4[7:6]);
    parallel_prefix mod100(temp_3[9:8], 2'b00, temp_4[9:8]);
    parallel_prefix mod101(temp_3[11:10], 2'b00, temp_4[11:10]);
    parallel_prefix mod102(temp_3[13:12], 2'b00, temp_4[13:12]);
    parallel_prefix mod103(temp_3[15:14], 2'b00, temp_4[15:14]);
    parallel_prefix mod104(temp_3[17:16], temp_4[15:14], temp_4[17:16]);
    parallel_prefix mod105(temp_3[19:18], temp_4[17:16], temp_4[19:18]);
    parallel_prefix mod106(temp_3[21:20], temp_4[19:18], temp_4[21:20]);
    parallel_prefix mod107(temp_3[23:22], temp_4[21:20], temp_4[23:22]);
    parallel_prefix mod108(temp_3[25:24], temp_4[23:22], temp_4[25:24]);
    parallel_prefix mod109(temp_3[27:26], temp_4[25:24], temp_4[27:26]);
    parallel_prefix mod110(temp_3[29:28], temp_4[27:26], temp_4[29:28]);
    parallel_prefix mod111(temp_3[31:30], temp_4[29:28], temp_4[31:30]);
    parallel_prefix mod112(temp_3[33:32], temp_4[31:30], temp_4[33:32]);
    parallel_prefix mod113(temp_3[35:34], temp_4[33:32], temp_4[35:34]);
    parallel_prefix mod114(temp_3[37:36], temp_4[35:34], temp_4[37:36]);
    parallel_prefix mod115(temp_3[39:38], temp_4[37:36], temp_4[39:38]);
    parallel_prefix mod116(temp_3[41:40], temp_4[39:38], temp_4[41:40]);
    parallel_prefix mod117(temp_3[43:42], temp_4[41:40], temp_4[43:42]);
    parallel_prefix mod118(temp_3[45:44], temp_4[43:42], temp_4[45:44]);
    parallel_prefix mod119(temp_3[47:46], temp_4[45:44], temp_4[47:46]);
    parallel_prefix mod120(temp_3[49:48], temp_4[47:46], temp_4[49:48]);
    parallel_prefix mod121(temp_3[51:50], temp_4[49:48], temp_4[51:50]);
    parallel_prefix mod122(temp_3[53:52], temp_4[51:50], temp_4[53:52]);
    parallel_prefix mod123(temp_3[55:54], temp_4[53:52], temp_4[55:54]);
    parallel_prefix mod124(temp_3[57:56], temp_4[55:54], temp_4[57:56]);
    parallel_prefix mod125(temp_3[59:58], temp_4[57:56], temp_4[59:58]);
    parallel_prefix mod126(temp_3[61:60], temp_4[59:58], temp_4[61:60]);
    parallel_prefix mod127(temp_3[63:62], temp_4[61:60], temp_4[63:62]);

endmodule
