module level_5 (
    input [63:0] temp_4, output [63:0] temp_5
);

    parallel_prefix mod128(temp_4[1:0], 2'b00, temp_5[1:0]);
    parallel_prefix mod129(temp_4[3:2], 2'b00, temp_5[3:2]);
    parallel_prefix mod130(temp_4[5:4], 2'b00, temp_5[5:4]);
    parallel_prefix mod131(temp_4[7:6], 2'b00, temp_5[7:6]);
    parallel_prefix mod132(temp_4[9:8], 2'b00, temp_5[9:8]);
    parallel_prefix mod133(temp_4[11:10], 2'b00, temp_5[11:10]);
    parallel_prefix mod134(temp_4[13:12], 2'b00, temp_5[13:12]);
    parallel_prefix mod135(temp_4[15:14], 2'b00, temp_5[15:14]);
    parallel_prefix mod136(temp_4[17:16], 2'b00, temp_5[17:16]);
    parallel_prefix mod137(temp_4[19:18], 2'b00, temp_5[19:18]);
    parallel_prefix mod138(temp_4[21:20], 2'b00, temp_5[21:20]);
    parallel_prefix mod139(temp_4[23:22], 2'b00, temp_5[23:22]);
    parallel_prefix mod140(temp_4[25:24], 2'b00, temp_5[25:24]);
    parallel_prefix mod141(temp_4[27:26], 2'b00, temp_5[27:26]);
    parallel_prefix mod142(temp_4[29:28], 2'b00, temp_5[29:28]);
    parallel_prefix mod143(temp_4[31:30], 2'b00, temp_5[31:30]);
    parallel_prefix mod144(temp_4[33:32], temp_5[31:30], temp_5[33:32]);
    parallel_prefix mod145(temp_4[35:34], temp_5[33:32], temp_5[35:34]);
    parallel_prefix mod146(temp_4[37:36], temp_5[35:34], temp_5[37:36]);
    parallel_prefix mod147(temp_4[39:38], temp_5[37:36], temp_5[39:38]);
    parallel_prefix mod148(temp_4[41:40], temp_5[39:38], temp_5[41:40]);
    parallel_prefix mod149(temp_4[43:42], temp_5[41:40], temp_5[43:42]);
    parallel_prefix mod150(temp_4[45:44], temp_5[43:42], temp_5[45:44]);
    parallel_prefix mod151(temp_4[47:46], temp_5[45:44], temp_5[47:46]);
    parallel_prefix mod152(temp_4[49:48], temp_5[47:46], temp_5[49:48]);
    parallel_prefix mod153(temp_4[51:50], temp_5[49:48], temp_5[51:50]);
    parallel_prefix mod154(temp_4[53:52], temp_5[51:50], temp_5[53:52]);
    parallel_prefix mod155(temp_4[55:54], temp_5[53:52], temp_5[55:54]);
    parallel_prefix mod156(temp_4[57:56], temp_5[55:54], temp_5[57:56]);
    parallel_prefix mod157(temp_4[59:58], temp_5[57:56], temp_5[59:58]);
    parallel_prefix mod158(temp_4[61:60], temp_5[59:58], temp_5[61:60]);
    parallel_prefix mod159(temp_4[63:62], temp_5[61:60], temp_5[63:62]);


endmodule
