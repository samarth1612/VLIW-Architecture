`include "include.v"

module processor ();
    
    RegisterFile rf ();
    
endmodule
