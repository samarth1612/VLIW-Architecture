`include "include.v"

module processor ();
    
    RegisterFile rf ();
    memory mem();
    
endmodule
