module level_2(
    input [63:0] temp_1, output [63:0] temp_2
);

    parallel_prefix mod32(temp_1[1:0], 2'b00, temp_2[1:0]);
    parallel_prefix mod33(temp_1[3:2], 2'b00, temp_2[3:2]);
    parallel_prefix mod34(temp_1[5:4], temp_2[3:2], temp_2[5:4]);
    parallel_prefix mod35(temp_1[7:6], temp_2[5:4], temp_2[7:6]);
    parallel_prefix mod36(temp_1[9:8], temp_2[7:6], temp_2[9:8]);
    parallel_prefix mod37(temp_1[11:10], temp_2[9:8], temp_2[11:10]);
    parallel_prefix mod38(temp_1[13:12], temp_2[11:10], temp_2[13:12]);
    parallel_prefix mod39(temp_1[15:14], temp_2[13:12], temp_2[15:14]);
    parallel_prefix mod40(temp_1[17:16], temp_2[15:14], temp_2[17:16]);
    parallel_prefix mod41(temp_1[19:18], temp_2[17:16], temp_2[19:18]);
    parallel_prefix mod42(temp_1[21:20], temp_2[19:18], temp_2[21:20]);
    parallel_prefix mod43(temp_1[23:22], temp_2[21:20], temp_2[23:22]);
    parallel_prefix mod44(temp_1[25:24], temp_2[23:22], temp_2[25:24]);
    parallel_prefix mod45(temp_1[27:26], temp_2[25:24], temp_2[27:26]);
    parallel_prefix mod46(temp_1[29:28], temp_2[27:26], temp_2[29:28]);
    parallel_prefix mod47(temp_1[31:30], temp_2[29:28], temp_2[31:30]);
    parallel_prefix mod48(temp_1[33:32], temp_2[31:30], temp_2[33:32]);
    parallel_prefix mod49(temp_1[35:34], temp_2[33:32], temp_2[35:34]);
    parallel_prefix mod50(temp_1[37:36], temp_2[35:34], temp_2[37:36]);
    parallel_prefix mod51(temp_1[39:38], temp_2[37:36], temp_2[39:38]);
    parallel_prefix mod52(temp_1[41:40], temp_2[39:38], temp_2[41:40]);
    parallel_prefix mod53(temp_1[43:42], temp_2[41:40], temp_2[43:42]);
    parallel_prefix mod54(temp_1[45:44], temp_2[43:42], temp_2[45:44]);
    parallel_prefix mod55(temp_1[47:46], temp_2[45:44], temp_2[47:46]);
    parallel_prefix mod56(temp_1[49:48], temp_2[47:46], temp_2[49:48]);
    parallel_prefix mod57(temp_1[51:50], temp_2[49:48], temp_2[51:50]);
    parallel_prefix mod58(temp_1[53:52], temp_2[51:50], temp_2[53:52]);
    parallel_prefix mod59(temp_1[55:54], temp_2[53:52], temp_2[55:54]);
    parallel_prefix mod60(temp_1[57:56], temp_2[55:54], temp_2[57:56]);
    parallel_prefix mod61(temp_1[59:58], temp_2[57:56], temp_2[59:58]);
    parallel_prefix mod62(temp_1[61:60], temp_2[59:58], temp_2[61:60]);
    parallel_prefix mod63(temp_1[63:62], temp_2[61:60], temp_2[63:62]);

endmodule
