module level_3(
    input [63:0] temp_2, output [63:0] temp_3
);

    parallel_prefix mod64(temp_2[1:0], 2'b00, temp_3[1:0]);
    parallel_prefix mod65(temp_2[3:2], 2'b00, temp_3[3:2]);
    parallel_prefix mod66(temp_2[5:4], 2'b00, temp_3[5:4]);
    parallel_prefix mod67(temp_2[7:6], 2'b00, temp_3[7:6]);
    parallel_prefix mod68(temp_2[9:8], temp_3[7:6], temp_3[9:8]);
    parallel_prefix mod69(temp_2[11:10], temp_3[9:8], temp_3[11:10]);
    parallel_prefix mod70(temp_2[13:12], temp_3[11:10], temp_3[13:12]);
    parallel_prefix mod71(temp_2[15:14], temp_3[13:12], temp_3[15:14]);
    parallel_prefix mod72(temp_2[17:16], temp_3[15:14], temp_3[17:16]);
    parallel_prefix mod73(temp_2[19:18], temp_3[17:16], temp_3[19:18]);
    parallel_prefix mod74(temp_2[21:20], temp_3[19:18], temp_3[21:20]);
    parallel_prefix mod75(temp_2[23:22], temp_3[21:20], temp_3[23:22]);
    parallel_prefix mod76(temp_2[25:24], temp_3[23:22], temp_3[25:24]);
    parallel_prefix mod77(temp_2[27:26], temp_3[25:24], temp_3[27:26]);
    parallel_prefix mod78(temp_2[29:28], temp_3[27:26], temp_3[29:28]);
    parallel_prefix mod79(temp_2[31:30], temp_3[29:28], temp_3[31:30]);
    parallel_prefix mod80(temp_2[33:32], temp_3[31:30], temp_3[33:32]);
    parallel_prefix mod81(temp_2[35:34], temp_3[33:32], temp_3[35:34]);
    parallel_prefix mod82(temp_2[37:36], temp_3[35:34], temp_3[37:36]);
    parallel_prefix mod83(temp_2[39:38], temp_3[37:36], temp_3[39:38]);
    parallel_prefix mod84(temp_2[41:40], temp_3[39:38], temp_3[41:40]);
    parallel_prefix mod85(temp_2[43:42], temp_3[41:40], temp_3[43:42]);
    parallel_prefix mod86(temp_2[45:44], temp_3[43:42], temp_3[45:44]);
    parallel_prefix mod87(temp_2[47:46], temp_3[45:44], temp_3[47:46]);
    parallel_prefix mod88(temp_2[49:48], temp_3[47:46], temp_3[49:48]);
    parallel_prefix mod89(temp_2[51:50], temp_3[49:48], temp_3[51:50]);
    parallel_prefix mod90(temp_2[53:52], temp_3[51:50], temp_3[53:52]);
    parallel_prefix mod91(temp_2[55:54], temp_3[53:52], temp_3[55:54]);
    parallel_prefix mod92(temp_2[57:56], temp_3[55:54], temp_3[57:56]);
    parallel_prefix mod93(temp_2[59:58], temp_3[57:56], temp_3[59:58]);
    parallel_prefix mod94(temp_2[61:60], temp_3[59:58], temp_3[61:60]);
    parallel_prefix mod95(temp_2[63:62], temp_3[61:60], temp_3[63:62]);

endmodule
